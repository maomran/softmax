`define DATALENGTH 32
module softmax(
		clk
		rst
		[`DATALENGTH-1:0] );